`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:34:50 11/18/2018 
// Design Name: 
// Module Name:    pack 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pack(
    input [1:0]a,
	 input [1:0]b,
	 input cin,
	 input [1:0]select,
	 output [3:0]out);
	alu

endmodule
